mux_add2 <= '';
mux_7sh <= '';
mux_a2 <= '';
mux_a3 <= "";
mux_d1 <= '';
mux_d2 <= '';
mux_op1 <= "";
mux_op2 <= "";
mux_dr <= '';
mux_rfd <= '';
mux_z2 <= '';
alu_op_sel <= '';
wr_mem <= '';
wr_rf <= '';
op1_check <= '';
op2_check <= '';
dest_cycle <= '';
source1_cycle <= "";
source2_cycle <= "";
mux_ao <= '';
valid_dest <= '';
lm_detected <= '';
sm_detected <= '';
